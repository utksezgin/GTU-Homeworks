module alu_ctrl(aluctrl, funcfield, aluop);

	input [5:0] aluop;
	input [6:0] funcfield;
	output [4:0] aluctrl; // add, addi
	
	
	
		
endmodule